// 8-3优先编码器
module lab2(
    input en,
    input[7:0] x,
    output[2:0] y,
    output i,
    output[6:0] hex
);
    assign i = en & (|x);
    wire[7:0] c;
    assign c[7] = x[7];
    assign c[6] = x[6] & (~x[7]);
    assign c[5] = x[5] & (~|x[7:6]);
    assign c[4] = x[4] & (~|x[7:5]);
    assign c[3] = x[3] & (~|x[7:4]);
    assign c[2] = x[2] & (~|x[7:3]);
    assign c[1] = x[1] & (~|x[7:2]);
    assign c[0] = x[0] & (~|x[7:1]);

    assign y = {3{en}} & ({3{c[0]}}&3'd0 | {3{c[1]}}&3'd1 | {3{c[2]}}&3'd2 | {3{c[3]}}&3'd3 | {3{c[4]}}&3'd4 | {3{c[5]}}&3'd5 | {3{c[6]}}&3'd6 | {3{c[7]}}&3'd7);

    assign hex = {7{en}} & (({7{y==3'd0}} &7'b1000000) | ({7{y==3'd1}} &7'b1111001) | ({7{y==3'd2}} &7'b0100100) | ({7{y==3'd3}} &7'b0110000) | ({7{y==3'd4}} &7'b0011001) | ({7{y==3'd5}} &7'b0010010) | ({7{y==3'd6}} &7'b0000010) | ({7{y==3'd7}} &7'b1111000));
endmodule

